
module uart_module (
	clk_clk,
	led_export,
	reset_reset_n,
	switch_export,
	uart_rxd,
	uart_txd,
	sdram_addr,
	sdram_ba,
	sdram_cas_n,
	sdram_cke,
	sdram_cs_n,
	sdram_dq,
	sdram_dqm,
	sdram_ras_n,
	sdram_we_n);	

	input		clk_clk;
	output	[7:0]	led_export;
	input		reset_reset_n;
	input	[7:0]	switch_export;
	input		uart_rxd;
	output		uart_txd;
	output	[11:0]	sdram_addr;
	output	[1:0]	sdram_ba;
	output		sdram_cas_n;
	output		sdram_cke;
	output		sdram_cs_n;
	inout	[15:0]	sdram_dq;
	output	[1:0]	sdram_dqm;
	output		sdram_ras_n;
	output		sdram_we_n;
endmodule
